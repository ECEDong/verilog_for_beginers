`define width 8
`define depth 8
`define addr  3